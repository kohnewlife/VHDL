library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY mips_control IS
	PORT(	opcode					:	IN	STD_LOGIC_VECTOR(5 DOWNTO 0);
			funct						:	IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			RegDst, ALUSrc			:	OUT STD_LOGIC;
			Jump, jal, Jr			:	OUT STD_LOGIC;
			Beq, Bne					:	OUT STD_LOGIC;
			MemRead, MemWrite		:	OUT STD_LOGIC;
			RegWrite, MemtoReg	:	OUT STD_LOGIC;
			ALUControl				:  OUT STD_LOGIC_VECTOR(3 DOWNTO 0)	);
END mips_control;

ARCHITECTURE Behavior OF mips_control IS

BEGIN 
	CASE opcode IS
		WHEN X"00" => 
			CASE funct IS
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
			END CASE;
		WHEN OTHERS => 
			CASE funct IS
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
				WHEN X"20" => 
					RegDst <= 
					ALUSrc <=
					Jump <=
					jal <=
					Jr <=
					Beq <=
					Bne <=
					MemRead <=
					MemWrite <=
					RegWrite <=
					MemtoReg <=
					ALUControl <=
			END CASE;
	END CASE;
			
END Behavior;